*2.8

r1 1 2 1
r2 2 3 2
c1 2 0 1u ic=0
v1 1 0 1
v2 3 0 2

.tran 10p 10u 0 uic
.control
run
set gnuplot_terminal=pdf/quit
gnuplot ../figs/2.8 v(2)
.endc

.end
